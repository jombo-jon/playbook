-------------------------------------------------------------------------------
-- Project name      : 
-- Project number    :
-- Customer          : 
--
-- Used Primitives   : 
--
-------------------------------------------------------------------------------
-- Description : 
-- 
-------------------------------------------------------------------------------

