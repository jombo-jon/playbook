-------------------------------------------------------------------------------
-- Project name      : {Project Name}
-- Project number    : {Project Number}
-- Customer          : {Customer} 
--
-- Used Primitives   : 
--
-------------------------------------------------------------------------------
-- Description : 
-- {Description} 
-------------------------------------------------------------------------------

