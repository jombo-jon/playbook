-------------------------------------------------------------------------------
-- Project name      : {Project Name}
-- Project number    : {Project Number}
-- Customer          : {CUstomer} 
--
-- Used Primitives   : 
--
-------------------------------------------------------------------------------
-- Description : 
-- 
-------------------------------------------------------------------------------
package FunctionPkg is

end FunctionPkg;

package body FunctionPkg is

end FunctionPkg;
