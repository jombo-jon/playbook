-- Test template VHD
