-- Package
