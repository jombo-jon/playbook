-------------------------------------------------------------------------------
-- Project name      : {Project Name}
-- Project number    : {Project Number}
-- Customer          : {Customer} 
--
-- Used Primitives   : 
--
-------------------------------------------------------------------------------
-- Description : 
-- 
-------------------------------------------------------------------------------
package {Package Name} is

  end {Package Name};

package body {Package Name} is

  end {Package Name};


